// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Booths_Multiplier
// --------------------------------------------------

module Booths_Multiplier (
    // Inputs
    // Outputs
);

endmodule
