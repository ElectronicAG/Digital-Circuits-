// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Multiplexer
// --------------------------------------------------

module Multiplexer (
    // Inputs
    // Outputs
);

endmodule
