// Date: 07/01/2026
// Autor: Alan Gomez
// Module: JK_Flip-Flop
// --------------------------------------------------

module JK_Flip-Flop (
    // Inputs
    // Outputs
);

endmodule
