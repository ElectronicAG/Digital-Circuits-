// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Moore_Sequence_Detector
// --------------------------------------------------

module Moore_Sequence_Detector (
    // Inputs
    // Outputs
);

endmodule
