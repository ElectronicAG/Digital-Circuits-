// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Priority_Encoder
// --------------------------------------------------

module Priority_Encoder (
    // Inputs
    // Outputs
);

endmodule
