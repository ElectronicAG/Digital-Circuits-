// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Synchronous_Counter
// --------------------------------------------------

module Synchronous_Counter (
    // Inputs
    // Outputs
);

endmodule
