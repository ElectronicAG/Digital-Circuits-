// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Demultiplexer
// --------------------------------------------------

module Demultiplexer (
    // Inputs
    // Outputs
);

endmodule
