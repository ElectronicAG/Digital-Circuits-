// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Comparator
// --------------------------------------------------

module Comparator (
    // Inputs
    // Outputs
);

endmodule
