// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Ripple_Carry_Adder
// --------------------------------------------------

module Ripple_Carry_Adder (
    // Inputs
    // Outputs
);

endmodule
