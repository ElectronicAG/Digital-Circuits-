// Date: 07/01/2026
// Autor: Alan Gomez
// Module: SR_Flip-Flop
// --------------------------------------------------

module SR_Flip-Flop (
    // Inputs
    // Outputs
);

endmodule
