// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Decoder
// --------------------------------------------------

module Decoder (
    // Inputs
    // Outputs
);

endmodule
