// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Encoder
// --------------------------------------------------

module Encoder (
    // Inputs
    // Outputs
);

endmodule
