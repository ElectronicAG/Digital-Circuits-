// Date: 07/01/2026
// Autor: Alan Gomez
// Module: 4-bit_Adder_Subtractor
// --------------------------------------------------

module 4-bit_Adder_Subtractor (
    // Inputs
    // Outputs
);

endmodule
