// Date: 07/01/2026
// Autor: Alan Gomez
// Module: Synchronous_FIFO
// --------------------------------------------------

module Synchronous_FIFO (
    // Inputs
    // Outputs
);

endmodule
